module Lab4(
);

endnoduke