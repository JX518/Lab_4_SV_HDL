//ALU should handle the calculations of 
	// next PC
	// addition
	// multiplication
	// comparison
	// nop
	// loading from mem

	// selecting immediate

module ALU(
	input logic [2:0] op,
	input logic [2:0] ra,
	input logic [2:0] rb,
	input logic [2:0] rd,   
	output logic [5:0] d	  
);
