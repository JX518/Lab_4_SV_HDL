module Lab4(	    
);
(* ram_init_file = "Lab4.mif" *) logic [11:0] mem[63:0];

assign *Instruction Code* = mem[*Program Counter*];

endmodule