//ALU should handle the calculations of 
	// next PC
	// addition
	// multiplication
	// comparison
	// nop
	// loading from mem

	// selecting immediate
